		--Decoder: address -> Chip Select 
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;

ENTITY CS_DEC IS
   PORT( 	
	address : IN  STD_LOGIC_VECTOR( 4  DOWNTO 0 );	-- ( A11 A5 A4 A3 A2 )
	CS		: OUT STD_LOGIC_VECTOR( 10 DOWNTO 0 )
	);
END CS_DEC;

ARCHITECTURE behavior OF CS_DEC IS				
BEGIN   
	WITH address SELECT
		CS <= "00000000001"  WHEN "10000", -- CS0 = 0x800 (LEDR)
			  "00000000010"  WHEN "10001", -- CS1 = 0x804 (HEX0) || 0x805 (HEX1)
			  "00000000100"  WHEN "10010", -- CS2 = 0x808 (HEX2) || 0x809 (HEX3)
			  "00000001000"  WHEN "10011", -- CS3 = 0x80C (HEX4) || 0x80D (HEX5)
			  "00000010000"  WHEN "10100", -- CS4 = 0x810 (SW)		
			  "00000100000"  WHEN "10101", -- CS5 = 0x814 (KEY)
			  "00001000000"  WHEN "10111", -- CS6 = 0x81C (BTCTL)
			  "00010000000"  WHEN "11000", -- CS6 = 0x820 (BTCNT)
			  "00100000000"  WHEN "11001", -- CS6 = 0x824 (BTCCR0)
			  "01000000000"  WHEN "11010", -- CS6 = 0x828 (BTCCR1)
			  "10000000000"  WHEN "11011", -- CS6 = 0x82C (IE) || 0x82D (IFG) || 0x82E (TYPE)
			  "00000000000"  WHEN others;
END behavior;


